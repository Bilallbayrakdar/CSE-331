library verilog;
use verilog.vl_types.all;
entity tb_main_control is
end tb_main_control;
