library verilog;
use verilog.vl_types.all;
entity tb_pc_handler is
end tb_pc_handler;
