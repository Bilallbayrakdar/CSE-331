library verilog;
use verilog.vl_types.all;
entity tb_mips32 is
end tb_mips32;
