library verilog;
use verilog.vl_types.all;
entity \tb_xor_\ is
end \tb_xor_\;
