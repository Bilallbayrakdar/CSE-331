module mips32_testbench();

endmodule