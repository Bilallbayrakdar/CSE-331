library verilog;
use verilog.vl_types.all;
entity tb_program_counter is
end tb_program_counter;
