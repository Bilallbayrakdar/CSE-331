library verilog;
use verilog.vl_types.all;
entity tb_r_type is
end tb_r_type;
