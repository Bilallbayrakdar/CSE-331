library verilog;
use verilog.vl_types.all;
entity tb_and32 is
end tb_and32;
