library verilog;
use verilog.vl_types.all;
entity adder_18_tb is
end adder_18_tb;
