library verilog;
use verilog.vl_types.all;
entity tb_is_zero is
end tb_is_zero;
