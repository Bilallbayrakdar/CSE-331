library verilog;
use verilog.vl_types.all;
entity tb_or32 is
end tb_or32;
