library verilog;
use verilog.vl_types.all;
entity tb_shifter_2 is
end tb_shifter_2;
