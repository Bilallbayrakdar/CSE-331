library verilog;
use verilog.vl_types.all;
entity tb_extender_16_32 is
end tb_extender_16_32;
