library verilog;
use verilog.vl_types.all;
entity tb_adder_32 is
end tb_adder_32;
