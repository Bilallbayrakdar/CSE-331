library verilog;
use verilog.vl_types.all;
entity tb_mips32_registers is
end tb_mips32_registers;
