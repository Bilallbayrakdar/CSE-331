library verilog;
use verilog.vl_types.all;
entity tb_alu_1 is
end tb_alu_1;
