library verilog;
use verilog.vl_types.all;
entity tb_alu_32 is
end tb_alu_32;
