library verilog;
use verilog.vl_types.all;
entity tb_zero_extender_32 is
end tb_zero_extender_32;
