library verilog;
use verilog.vl_types.all;
entity tb_mux_4_1 is
end tb_mux_4_1;
