library verilog;
use verilog.vl_types.all;
entity tb_comparator_32 is
end tb_comparator_32;
