library verilog;
use verilog.vl_types.all;
entity tb_32_mux_2_1 is
end tb_32_mux_2_1;
